module demux_tb;

